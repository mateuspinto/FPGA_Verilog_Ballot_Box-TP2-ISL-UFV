module bcd7convert(bcd, SeteSegmentos, clock);

    output reg [6:0] SeteSegmentos;

    input[3:0] bcd;
    input clock;

    always @(posedge clock) begin

        case(bcd)

            4'b0000: SeteSegmentos = 7'b1000000;
            4'b0001: SeteSegmentos = 7'b1111001;
            4'b0010: SeteSegmentos = 7'b0100100;
            4'b0011: SeteSegmentos = 7'b0110000;
            4'b0100: SeteSegmentos = 7'b0011001;
            4'b0101: SeteSegmentos = 7'b0010010;
            4'b0110: SeteSegmentos = 7'b0000010;
            4'b0111: SeteSegmentos = 7'b1111000;
            4'b1000: SeteSegmentos = 7'b0000000;
            4'b1001: SeteSegmentos = 7'b0010000;
            4'b1010: SeteSegmentos = 7'b1111111;
            4'b1011: SeteSegmentos = 7'b1000110;
				4'b1100: SeteSegmentos = 7'b0101011;

        endcase

    end

endmodule